module (ip_0,ip_1,ip_2,ip_3,ip_4,ip_5,ip_6,ip_7,ip_8,ip_9,ip_10,ip_11,ip_12,ip_13,ip_14,ip_15,ip_16,ip_17,ip_18,ip_19,ip_20,ip_21,ip_22,ip_23,ip_24,ip_25,ip_26,ip_27,ip_28,ip_29,ip_30,ip_31,ip_32,ip_33,ip_34,ip_35,ip_36,ip_37,ip_38,ip_39,ip_40,ip_41,ip_42,ip_43,ip_44,ip_45,ip_46,ip_47,ip_48,ip_49,ip_50,ip_51,ip_52,ip_53,ip_54,ip_55,ip_56,ip_57,ip_58,ip_59,ip_60,ip_61,ip_62,ip_63, o1);
input ip_0, ip_1, ip_2, ip_3, ip_4, ip_5, ip_6, ip_7, ip_8, ip_9, ip_10, ip_11, ip_12, ip_13, ip_14, ip_15, ip_16, ip_17, ip_18, ip_19, ip_20, ip_21, ip_22, ip_23, ip_24, ip_25, ip_26, ip_27, ip_28, ip_29, ip_30, ip_31, ip_32, ip_33, ip_34, ip_35, ip_36, ip_37, ip_38, ip_39, ip_40, ip_41, ip_42, ip_43, ip_44, ip_45, ip_46, ip_47, ip_48, ip_49, ip_50, ip_51, ip_52, ip_53, ip_54, ip_55, ip_56, ip_57, ip_58, ip_59, ip_60, ip_61, ip_62, ip_63;
output o1;
wire w_0;

assign o1 = ip_0;
endmodule
